<svg id="Layer_1" data-name="Layer 1" xmlns="http://www.w3.org/2000/svg" viewBox="0 0 48 48"><defs><style>.cls-1{fill:none;stroke:#054d7f;stroke-linecap:round;stroke-miterlimit:10;stroke-width:0.574px;}.cls-2{fill:#fff;}</style></defs><title>Single bed</title><path class="cls-1" d="M37.689,21.168V11.223a2.308,2.308,0,0,0-2.308-2.308H12.541a2.308,2.308,0,0,0-2.308,2.308v9.945"/><path class="cls-1" d="M17.924,23.115v-5.64A1.879,1.879,0,0,1,19.8,15.6H28.2a1.879,1.879,0,0,1,1.88,1.879v5.64"/><path class="cls-1" d="M40.011,29.507v9.578H34.774v-2.82a2.417,2.417,0,0,0-2.417-2.417H15.643a2.417,2.417,0,0,0-2.417,2.417v2.82H7.989V25.331a2.216,2.216,0,0,1,2.216-2.216H37.8a2.216,2.216,0,0,1,2.216,2.216Z"/><path class="cls-2" d="M24,27.094a34.425,34.425,0,0,1,14.355,2.812V25.331a.56.56,0,0,0-.559-.56H10.205a.56.56,0,0,0-.56.56v4.575A34.425,34.425,0,0,1,24,27.094Z"/></svg>